# ====================================================================
#
#	opencores_ethmac_eth_drivers.cdl
#
#	OpenCores ETHMAC ethernet driver
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2003, 2004 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Piotr Skrzypek
# Original data:
# Contributors:
# Date:           2012-04-10
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_ETH_OPENCORES_ETHMAC {

    display       "OpenCores ETHMAC ethernet driver"
    description   "Ethernet driver for OpenCores ETHMAC controller."

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if     CYGPKG_IO_ETH_DRIVERS

    implements    CYGHWR_NET_DRIVERS
    implements    CYGHWR_NET_DRIVER_ETH0

    compile       -library=libextras.a if_ethmac.c

    cdl_option CYGPKG_DEVS_ETH_OPENCORES_ETHMAC_MACADDR {
        display "Ethernet station (MAC) address for eth0"
        flavor  data
        default_value {"0x12, 0x34, 0x56, 0x78, 0x9A, 0xBC"}
        description   "The default ethernet station address. This is the
                       MAC address used when no value is found in the
                       RedBoot FLASH configuration field."
    }

    cdl_option CYGPKG_DEVS_ETH_OPENCORES_ETHMAC_INT {
        display "Interrupt vector number"
        flavor  data
        default_value { 4 }
        description   "
            This is the number of PIC channel that ETHMAC is connected
            to."
    }

    cdl_option CYGPKG_DEVS_ETH_OPENCORES_ETHMAC_INT_PRIO {
        display "Interrupt priority"
        flavor  data
        default_value { 4 }
        description   "
            Priority of delayed interrupt routine that takes care
            of ETHMAC."
    }

    cdl_option CYGPKG_DEVS_ETH_OPENCORES_ETHMAC_TXBUF_COUNT {
        display "Number of transmit buffers"
        flavor  data
        default_value { 1 }
        legal_values 1 to 64
        description   "
            The number of transmit buffers. More buffers help
            increse the throughput, but require maintenance time
            and  memory."
    }

    cdl_option CYGPKG_DEVS_ETH_OPENCORES_ETHMAC_RXBUF_COUNT {
        display "Number of receive buffers"
        flavor  data
        default_value { 1 }
        legal_values 1 to 64
        description   "
            The number of receive buffers. More buffers prevent
            missing packets, but require more maintenance time
            and memory."
    }

    cdl_option CYGPKG_DEVS_ETH_OPENCORES_ETHMAC_PACKETLEN {
        display "Maximum frame length"
        flavor  data
        default_value { 1536 }
        description   "
            Specify maximum packet length. This value will be
            programmed into the MAC. It is also a size of receive
            buffers."
    }

    cdl_option CYGPKG_DEVS_ETH_OPENCORES_ETHMAC_FULLDUPLEX {
        display "Enable full duplex transmission"
        flavor  bool
        default_value { 1 }
        description   "
            Enable full duplex when configuring ETHMAC."
    }

    cdl_component CYGPKG_DEVS_ETH_OPENCORES_ETHMAC_OPTIONS {
        display "ETHMAC controller driver build options"
        flavor  none
        no_define

        cdl_option CYGPKG_DEVS_ETH_OPENCORES_ETHMAC_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS" }
            description   "
                This option modifies the set of compiler flags for
                building the ETHMAC controller driver package.
                These flags are used in addition to the set of global
                flags."
        }
    }


}
# EOF opencores_ethmac_eth_drivers.cdl
