# ====================================================================
#
#      hal_openrisc.cdl
#
#      OpenRISC architectural HAL package configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2003 Free Software Foundation, Inc.                        
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      sfurman
# Original data:  bartv, nickg
# Contributors:   jskov
# Date:           2003-02-28
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_OPENRISC {
    display "OpenRISC architecture"
    parent        CYGPKG_HAL
    hardware
    include_dir   cyg/hal
    define_header hal_openrisc.h
    description   "
        The OpenRISC architecture HAL package provides generic support
        for this processor architecture. It is also necessary to
        select a specific target platform HAL package."

    compile       context.S vectors.S hal_misc.c openrisc_stub.c

    implements    CYGINT_HAL_DEBUG_GDB_STUBS
    implements    CYGINT_HAL_DEBUG_GDB_STUBS_BREAK

    make {
        <PREFIX>/lib/vectors.o : <PACKAGE>/src/vectors.S
        $(CC) -Wp,-MD,vectors.tmp $(INCLUDE_PATH) $(CFLAGS) -c -o $@ $<
        @echo $@ ": \\" > $(notdir $@).deps
        @tail -n +2 vectors.tmp >> $(notdir $@).deps
        @echo >> $(notdir $@).deps
        @rm vectors.tmp
    }

    define_proc {
        puts $::cdl_header "#define HAL_ARCH_PROGRAM_NEW_STACK hal_arch_program_new_stack"
    }

    cdl_option CYGBLD_LINKER_SCRIPT {
        display "Linker script"
        flavor data
        no_define
        calculated  { "src/openrisc.ld" }
    }

    make {
        <PREFIX>/lib/target.ld: <PACKAGE>/src/openrisc.ld
        $(CC) -E -P -Wp,-MD,target.tmp -DEXTRAS=1 -xc $(INCLUDE_PATH) $(ACTUAL_CFLAGS) -o $@ $<
        @echo $@ ": \\" > $(notdir $@).deps
        @tail -n +2 target.tmp >> $(notdir $@).deps
        @echo >> $(notdir $@).deps
        @rm target.tmp
    }

    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        legal_values  {"RAM" "ROM" "JTAG"}
        default_value {"JTAG"}
        no_define
        define -file system.h CYG_HAL_STARTUP
        description   "
            Selects whether code initially runs from ROM or RAM.  In the case of ROM startup,
            it's possible for the code to be copied into RAM and executed there."
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { CYG_HAL_STARTUP == "ROM" ? "openrisc_orpsoc_rom" : \
                                                "openrisc_orpsoc_ram" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { CYG_HAL_STARTUP == "ROM" ? "<pkgconf/mlt_openrisc_orpsoc_rom.ldi>" : \
                                                    "<pkgconf/mlt_openrisc_orpsoc_ram.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { CYG_HAL_STARTUP == "ROM" ? "<pkgconf/mlt_openrisc_orpsoc_rom.h>" : \
                                                    "<pkgconf/mlt_openrisc_orpsoc_ram.h>" }
        }
    }

    # Real-time clock/counter specifics
    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants."
        flavor        none

        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            default_value 1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            default_value 100
        }
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
            default_value {CYGHWR_HAL_OPENRISC_CPU_FREQ * 1000000 / CYGNUM_HAL_RTC_DENOMINATOR}
            description   "
                The tick timer facility is used
                to drive the eCos kernel RTC. The count register
                increments at the CPU clock speed.  By default, 100 Hz"
        }
    }

    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        description   "
            Global build options including control over
            compiler flags, linker flags and choice of toolchain."


        parent  CYGPKG_NONE

        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "or32-elf" }
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { CYGBLD_GLOBAL_WARNFLAGS . 
                            "-g -O2 -fno-omit-frame-pointer -fno-rtti -fno-exceptions " . 
                            (CYGHWR_MUL_IMPLEMENTED ? "-mhard-mul " : "-msoft-mul ") .
                            (CYGHWR_DIV_IMPLEMENTED ? "-mhard-div " : "-msoft-div ") .
                            (CYGHWR_FPU_IMPLEMENTED ? "-mhard-float " : "-msoft-float ") }
            description   "
                This option controls the global compiler flags which
                are used to compile all packages by
                default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { "-g -O2 -nostdlib -Wl,--gc-sections -Wl,-static " . 
                            (CYGHWR_MUL_IMPLEMENTED ? "-mhard-mul " : "-msoft-mul ") .
                            (CYGHWR_DIV_IMPLEMENTED ? "-mhard-div " : "-msoft-div ") .
                            (CYGHWR_FPU_IMPLEMENTED ? "-mhard-float " : "-msoft-float ") }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }
    }

    cdl_option CYGBLD_BUILD_GDB_STUBS {
        display "Build GDB stub ROM image"
        default_value 0
        parent CYGBLD_GLOBAL_OPTIONS
        requires { CYG_HAL_STARTUP == "ROM" }
        requires CYGSEM_HAL_ROM_MONITOR
        requires CYGBLD_BUILD_COMMON_GDB_STUBS
        requires CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
        requires ! CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT
        requires ! CYGDBG_HAL_DEBUG_GDB_THREAD_SUPPORT
        requires ! CYGDBG_HAL_COMMON_INTERRUPTS_SAVE_MINIMUM_CONTEXT
        requires ! CYGDBG_HAL_COMMON_CONTEXT_SAVE_MINIMUM
        no_define
        description "
                This option enables the building of the GDB stubs for the
                board. The common HAL controls takes care of most of the
                build process, but the final conversion from ELF image to
                binary data is handled by the platform CDL, allowing
                relocation of the data if necessary."

        make -priority 320 {
            <PREFIX>/bin/gdb_module.bin : <PREFIX>/bin/gdb_module.img
            $(OBJCOPY) -O binary $< $@
        }
    }

    cdl_option CYGNUM_HAL_BREAKPOINT_LIST_SIZE {
        display       "Number of breakpoints supported by the HAL."
        flavor        data
        default_value 25
        description   "
            This option determines the number of breakpoints supported by the HAL."
    }

    cdl_option CYGSEM_HAL_USE_ROM_MONITOR {
        display       "Work with a ROM monitor"
        flavor        bool
        default_value { CYG_HAL_STARTUP == "RAM" ? 1 : 0 }
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "RAM" }
        description   "
            Allow coexistence with ROM monitor (CygMon or GDB stubs) by
            only initializing interrupt vectors on startup, thus leaving
            exception handling to the ROM monitor."
    }

    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 0
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "ROM" }
        description   "
            Enable this option if this program is to be used as a ROM monitor,
            i.e. applications will be loaded into RAM on the board, and this
            ROM monitor may process exceptions or interrupts generated from the
            application. This enables features such as utilizing a separate
            interrupt stack when exceptions are generated."
    }

    cdl_component CYGPKG_REDBOOT_HAL_OPTIONS {
        display       "Redboot HAL options"
        flavor        none
        no_define
        parent        CYGPKG_REDBOOT
        active_if     CYGPKG_REDBOOT
        description   "
            This option lists the target's requirements for a valid Redboot
            configuration."

        cdl_option CYGBLD_BUILD_REDBOOT_BIN {
            display       "Build Redboot ROM binary image"
            active_if     CYGBLD_BUILD_REDBOOT
            default_value 1
            no_define
            description "This option enables the conversion of the Redboot ELF
                         image to a binary image suitable for ROM programming."

            compile -library=libextras.a

            make -priority 325 {
                <PREFIX>/bin/redboot.srec : <PREFIX>/bin/redboot.elf
                $(OBJCOPY) --strip-all $< $(@:.srec=.img)
                $(OBJCOPY) -O srec $< $@
            }
        }
    }

    cdl_option CYGHWR_HAL_OPENRISC_CPU_FREQ {
        display "CPU frequency"
        flavor  data
        legal_values 0 to 1000000
        default_value 50
        description "
           This option contains the frequency of the CPU in MegaHertz.
           Choose the frequency to match the processor you have. This
           may affect thing like serial device, interval clock and
           memory access speed settings."
    }

    cdl_option CYGHWR_MUL_IMPLEMENTED {
        display       "Hardware multiplier implemented"
        flavor        bool
        default_value 1
        description   "
            Select this option only if hardware multiplier is
            implemented."
    }

    cdl_option CYGHWR_DIV_IMPLEMENTED {
        display       "Hardware divisor implemented"
        flavor        bool
        default_value 1
        description   "
            Select this option only if hardware division is
            implemented."
    }

    cdl_option CYGHWR_FPU_IMPLEMENTED {
        display       "Hardware FPU implemented"
        flavor        bool
        default_value 0
        description   "
            Select this option only if FPU is implemented."
    }

    cdl_component CYGHWR_CACHE {

        display "Cache"
        flavor none
        description "
           Cache is optional in the OpenRISC architecture. Removing 
           cache is a common way to save hardware space."

        cdl_option CYGHWR_ICACHE_IMPLEMENTED {
            display       "Instruction cache implemented"
            flavor        bool
            default_value 1
            description   "
                Select this option only if instruction cache is 
                implemented."
        }

        cdl_option CYGHWR_ICACHE_SIZE {
            display       "Instruction cache size"
            active_if     CYGHWR_ICACHE_IMPLEMENTED
            flavor        data
            legal_values  4096 8192
            default_value 8192
            description   "
                Size of the instruction cache."
        }

        cdl_option CYGHWR_DCACHE_IMPLEMENTED {
            display       "Data cache implemented"
            flavor        bool
            default_value 1
            description   "
                Select this option only if data cache is 
                implemented."
        }

        cdl_option CYGHWR_DCACHE_SIZE {
            display       "Data cache size"
            active_if     CYGHWR_DCACHE_IMPLEMENTED
            flavor        data
            legal_values  4096 8192
            default_value 4096
            description   "
                Size of the data cache."
        }

    }

}

# EOF hal_openrisc.cdl
