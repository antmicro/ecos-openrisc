cdl_package CYGPKG_DEVS_SERIAL_OPENCORES_16550 {
    display         "OpenCores 16550 driver implementation"

    parent        CYGPKG_IO_SERIAL_DEVICES
    active_if     CYGPKG_IO_SERIAL


    requires      CYGPKG_ERROR
    include_dir     cyg/io
    description   "
        Enables serial device drivers for openrisc."


    # FIXME: This really belongs in the GENERIC_16X5X package
    cdl_interface CYGINT_IO_SERIAL_GENERIC_16X5X_REQUIRED {
        display   "Generic 16x5x serial driver required"
    }

    define_proc {
        puts $::cdl_system_header "/***** serial driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_GENERIC_16X5X_INL <cyg/io/opencores_16550_ser.inl>"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_GENERIC_16X5X_CFG <pkgconf/devs_serial_opencores_16550.h>"
        puts $::cdl_system_header "/*****  serial driver proc output end  *****/"
    }

cdl_component CYGPKG_IO_SERIAL_OPENCORES_SERIAL0 {
    display       "Serial port 0 driver"
    flavor        bool
    default_value 1
    description   "
        This option includes the serial device driver for port 0"


    implements    CYGINT_IO_SERIAL_GENERIC_16X5X_REQUIRED


    cdl_option CYGDAT_IO_SERIAL_OPENCORES_SERIAL0_NAME {
        display       "Device name"
        flavor        data
        default_value {"\"/dev/ser0\""}
        description   "
            This option specifies the device name port."
    }

    cdl_option CYGNUM_IO_SERIAL_OPENCORES_SERIAL0_BAUD {
        display       "Baud rate"
        flavor        data
        legal_values  { 1200 1800 2400 3600 4800 7200 9600
                        14400 19200 38400 57600 115200
        }
        default_value 115200
        description   "
            This option specifies the default baud rate (speed)"
    }

    cdl_option CYGNUM_IO_SERIAL_OPENCORES_SERIAL0_BUFSIZE {
        display       "Buffer size"
        flavor        data
        legal_values  0 to 8192
        default_value 128
        description   "
            This option specifies the size of the internal buffers used"
    }

    cdl_option CYGNUM_IO_SERIAL_OPENCORES_SERIAL0_IOBASE {
        display "I/O base address for the serial port "
        flavor    data
        legal_values 0 to 0xFFFFFFE0
        default_value 0x90000000
        description "
        This option specifies the I/O address"
    }

    cdl_option CYGNUM_IO_SERIAL_OPENCORES_SERIAL0_INT {
        display "INT for the serial port 0"
        flavor    data
        legal_values 2 to 21
        default_value 2
        description "
        This option specifies the interrupt vector for serial port 0."
   }
}
    cdl_component CYGPKG_IO_SERIAL_OPENCORES_TESTING {
        display    "Testing parameters"
        flavor     bool
        calculated 1
        active_if  CYGPKG_DEVS_SERIAL_OPENCORES_16550

        cdl_option CYGPRI_SER_TEST_SER_DEV {
            display       "Serial device used for testing"
            flavor        data
            default_value { CYGDAT_IO_SERIAL_OPENCORES_SERIAL0_NAME }
        }

        define_proc {
            puts $::cdl_header "#define CYGPRI_SER_TEST_CRASH_ID \"opencores\""
            puts $::cdl_header "#define CYGPRI_SER_TEST_TTY_DEV  \"/dev/tty0\""
        }
    }

}
