##=============================================================================
##
##      spi_simple_spi.cdl
##
##      OpenCores simple_spi driver configuration options.
##
##=============================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2008, 2009, 2011 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
##=============================================================================
#######DESCRIPTIONBEGIN####
##
## Author(s):   Piotr Skrzypek
## Date:        2012-05-14
##
######DESCRIPTIONEND####
##
##=============================================================================

cdl_package CYGPKG_DEVS_SPI_OPENCORES_SIMPLE_SPI {

    display       "OpenCores simple_spi driver"

    include_dir   cyg/io

    parent        CYGPKG_IO_SPI
    active_if     CYGPKG_IO_SPI

    compile       spi_simple_spi.c

    description   "
        This package provides SPI driver support for simple_spi project
        hosted on OpenCores."

    cdl_option CYGNUM_DEVS_SPI_OPENCORES_SIMPLE_SPI_COUNT {
        display       "Number of busses"
        flavor        data
        default_value 1
        description   "Enter the number of SPI busses in SoC."
    }

    cdl_option CYGNUM_DEVS_SPI_OPENCORES_SIMPLE_SPI_INT_PRI {
        display       "Interrupt priority"
        flavor        data
        default_value 5
    }

    cdl_option CYGNUM_DEVS_SPI_OPENCORES_SIMPLE_SPI_INTS {
        display       "Interrupt vectors"
        flavor        data
        default_value 6
        description   "Provide a comma separated list of interrupt vectors
                       connected to each bus."
    }

    cdl_option CYGNUM_DEVS_SPI_OPENCORES_SIMPLE_SPI_BUS_SPEED {
        display       "Bus speed"
        flavor        data
        default_value 50
        description   "Enter the speed of the bus that SPI is connected to.
                       Speed is in MHz. Needed to determine prescalers for
                       given device speeds."
    }

}
# EOF spi_simple_spi.cdl
