# ====================================================================
#
#      devs_disk_opencores_sdcmsc.cdl
#
#      Support for SDCard Mass Storage Controller
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2004, 2005, 2006 Free Software Foundation, Inc.            
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Piotr Skrzypek
# Date:           2012-05-01
#
#####DESCRIPTIONEND####
# ====================================================================

cdl_package CYGPKG_DEVS_DISK_OPENCORES_SDCMSC {
    display     "Disk driver for SDCard Mass Storage Controller"

    include_dir cyg/io
    
    parent      CYGPKG_IO_DISK_DEVICES
    active_if   CYGPKG_IO_DISK

    compile     -library=libextras.a if_sdcmsc.c
    requires    CYGPKG_ERROR CYGPKG_LIBC_STRING 

    description "
        This is a disk driver for SD Card Mass Storage Controller
        peripheral available at openCores."
	
    cdl_option CYGDAT_DEVS_DISK_OPENCORES_SDCMSC_DISK0_NAME {
        display		"Device name for the MMC/SPI disk 0 device"
        flavor		data
        default_value	{ "\"/dev/mmcdisk0/\"" }
        description "
            This is the device name used to access the raw disk device
            in eCos, for example for mount operations. Note that the
            trailing slash must be present."
        }
	
}

# EOF devs_disk_opencores_sdcmsc.cdl
